interface Sys_IF;
    logic clk_user;
    logic clk_hmc;  
    logic res_n_user; 
    logic res_n_hmc;
endinterface :Sys_IF
