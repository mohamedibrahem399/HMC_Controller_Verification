
package AXI_Req_pckg;
   import uvm_pkg::*;
`include "uvm_macros.svh"
 
   
  `include "CMD_DATA_TYPES.svh"
  `include "AXI_Req_Sequence_Item.svh"
  `include "Sequence.svh"
  `include "AXI_Sequencer.svh"
  `include "AXI_Req_Driver.svh"
  `include "AXI_Req_Monitor.svh"
  `include "AXI_Req_Agent.svh"
  `include "AXI_Req_Scoreboard.svh"
  `include "AXI_Req_Env.svh"
 
endpackage : AXI_Req_pckg
